    Mac OS X            	   2  >     p                                      ATTR      p   �   �                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl     4   <  com.apple.quarantine xse_    e �0     }i8Q�A��'���oL                                                      q/0081;5efc5eb1;Chrome;03B7D014-5A3B-4F62-867F-91E5F84FCE3C 